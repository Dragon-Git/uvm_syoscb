//----------------------------------------------------------------------
//   Copyright 2005-2022 SyoSil ApS
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------
  ////////////////////////////////////////////////////////////////////////////
  // TB Parameters
  ////////////////////////////////////////////////////////////////////////////

  // Number of scoreboards for scb_env
  localparam int unsigned NO_OF_SCB               = 2;

  // Number of scoreboards for scbs env
  localparam int unsigned NO_OF_SCBS              = 10;
